library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity principal is
    Port ( CLK  : in STD_LOGIC;                           -- Entrada de reloj
           SIN  : in STD_LOGIC;                           -- Entrada de datos
			  PULSADOR : in STD_LOGIC;                       -- Entrada Pulsador HORA/FECHA
			  LEDS : out STD_LOGIC_VECTOR (6 downto 0);      -- Salida LEDS d�a de la semana
           AN   : out STD_LOGIC_VECTOR (3 downto 0);      -- Control de displays
           SEG7 : out STD_LOGIC_VECTOR (6 downto 0));     -- Segmentos de displays
end principal;

architecture a_principal of principal is

-- Constantes del circuito (umbrales de decisi�n)

constant UMBRAL1 : STD_LOGIC_VECTOR (5 downto 0) := "100010"; -- 34 (Umbral comparador 1)
constant UMBRAL2 : STD_LOGIC_VECTOR (5 downto 0) := "100110"; -- 38 (Umbral comparador 2)

signal CLK_OUT : STD_LOGIC;        -- Se�al utilizada para las entradas que precisan la se�al CLK_M de 40 Hz
signal NQ0 : STD_LOGIC_VECTOR (39 downto 0);  -- Se�al que comunica la salida del registro de desplazamiento de 40 bits con el sumador.
signal NQ1 : STD_LOGIC_VECTOR (5 downto 0);   -- Se�al que comnica la salida del sumador con las entradas de los dos comparadores.
signal PGTQ1 : STD_LOGIC;                     -- Salida P>Q del comparador 1, corresponde a la primera entrada de la puerta AND.
signal PLEQ1 : STD_LOGIC;                     -- Salida P<=Q del comparador 1, corresponde a la segunda condici�n del aut�mata (SUM = U1).
signal PGTQ2 : STD_LOGIC;                     -- Salida P>Q del comparador 2.
signal PLEQ2 : STD_LOGIC;                     -- Salida P<=Q del comparador 2, corresponde a la segunda entrada de la puerta AND.
signal NQ2 : STD_LOGIC;                       -- Salida de la puerta AND, corresponde a la primera condici�n del aut�mata(U1 < SUM = U2).
signal NQ3 : STD_LOGIC;                       -- Salida del aut�mata, corresponde al Dato a cargar en el registro de desplazamiento de 14 bits.
signal NQ4 : STD_LOGIC;                       -- Salida del aut�mata, corresponde al ENABLE del registro de desplazamiento de 14 bits.
signal NQ5 : STD_LOGIC;                       -- Salida del aut�mata, corresponde al ENABLE del registro de validaci�n.
signal NQ6 : STD_LOGIC_VECTOR (30 downto 0);  -- Salida del registro de desplazamiento de 14 bits y entrada del registro de validaci�n.
signal NQ7 : STD_LOGIC_VECTOR (30 downto 0);  -- Salida del registro de validaci�n y entrada del m�dulo de visualizaci�n.
 

component gen_reloj
   Port ( CLK : in STD_LOGIC;         -- Reloj de la FPGA
          CLK_M : out STD_LOGIC);     -- Reloj de frecuencia dividida

end component;

component reg_desp40
   Port ( SIN : in STD_LOGIC;                          -- Datos de entrada serie
          CLK : in STD_LOGIC;                          -- Reloj de muestreo
          Q : out STD_LOGIC_VECTOR (39 downto 0));     -- Salida paralelo

end component;

component sumador40
   Port ( ENT : in STD_LOGIC_VECTOR (39 downto 0);
          SAL : out STD_LOGIC_VECTOR (5 downto 0));

end component;

component comparador
   Port ( P : in STD_LOGIC_VECTOR (5 downto 0);
          Q : in STD_LOGIC_VECTOR (5 downto 0);
          PGTQ : out STD_LOGIC;
          PLEQ : out STD_LOGIC);

end component;

component AND_2
   Port ( A : in STD_LOGIC;
          B : in STD_LOGIC;
          S : out STD_LOGIC);

end component;

component reg_desp
   Port ( SIN : in STD_LOGIC;                             -- Datos de entrada serie
          CLK : in STD_LOGIC;                             -- Reloj CLK_M
          EN : in STD_LOGIC;                              -- Enable
          Q : out STD_LOGIC_VECTOR (30 downto 0));        -- Salida paralelo

end component;
component registro
   Port ( ENTRADA : in STD_LOGIC_VECTOR (30 downto 0);
          SALIDA : out STD_LOGIC_VECTOR (30 downto 0);
          EN : in STD_LOGIC;                                   -- Enable
          RCLK : in STD_LOGIC);

end component;

component automata
   Port ( CLK : in STD_LOGIC;             -- Reloj del aut�mata
          C0 : in STD_LOGIC;              -- Condici�n de decision para "0"
          C1 : in STD_LOGIC;              -- Condici�n de decisi�n para "1"
          DATO : out STD_LOGIC;           -- Datos a cargar
          CAPTUR : out STD_LOGIC;         -- Enable del reg. de desplaz.
          VALID : out STD_LOGIC);         -- Activaci�n registro

end component;

component visualizacion
   Port ( E0 : in STD_LOGIC_VECTOR (3 downto 0);       -- Entrada MUX 0
          E1 : in STD_LOGIC_VECTOR (3 downto 0);       -- Entrada MUX 1
          E2 : in STD_LOGIC_VECTOR (3 downto 0);       -- Entrada MUX 2
          E3 : in STD_LOGIC_VECTOR (3 downto 0);       -- Entrada MUX 3
          E4 : in STD_LOGIC_VECTOR (3 downto 0);       -- Entrada MUX 4.
          E5 : in STD_LOGIC_VECTOR (3 downto 0);       -- Entrada MUX 5.
          E6 : in STD_LOGIC_VECTOR (3 downto 0);       -- Entrada MUX 6.
          E7 : in STD_LOGIC_VECTOR (3 downto 0);       -- Entrada MUX 7.
			 E8 : in STD_LOGIC_VECTOR (2 downto 0);       -- Entrada bits D�a semana.   
			 PULSADOR : in STD_LOGIC;                     -- Pulsador HORA/FECHA
			 CLK : in STD_LOGIC;                          -- Entrada de reloj FPGA
			 LEDS : out STD_LOGIC_VECTOR ( 6 downto 0);   -- LEDS salida d�a semana
          SEG7 : out STD_LOGIC_VECTOR (6 downto 0);    -- Salida para los displays
          AN : out STD_LOGIC_VECTOR (3 downto 0));     -- Activaci�n individual

end component;

begin

U1 : gen_reloj  -- Generador de reloj
       port map (
		   CLK => CLK,
			CLK_M => CLK_OUT
			);
			
U2 : reg_desp40  -- Registro de desplazamiento de 40 bits
       port map (
		   SIN => SIN,
			CLK => CLK_OUT,
			Q => NQ0
			);
			
U3 : sumador40  -- Integrador (sumador)
       port map (
         ENT => NQ0,
         SAL => NQ1
         );			
			
U4 : comparador -- Comparador 1
       port map (
		   P => NQ1,
			Q => UMBRAL1,
			PGTQ => PGTQ1,
			PLEQ => PLEQ1
			);
			
U5 : comparador -- Comparador 2
       port map (
		   P => NQ1,
			Q => UMBRAL2,
			PGTQ => PGTQ2,
			PLEQ => PLEQ2
			);
			
U6 : AND_2 -- Puerta AND
       port map (
		   A => PGTQ1,
			B => PLEQ2,
			S => NQ2
			);
			
U7 : automata -- Automata de MOORE
       port map (
		   CLK => CLK_OUT,
			C0 => NQ2,
			C1 => PLEQ1,
			DATO => NQ3,
			CAPTUR => NQ4,
			VALID => NQ5
			);
			
U8 : reg_desp  -- Registro de desplazamiento
       port map (
		   SIN => NQ3,
		   CLK => CLK_OUT,
		   EN => NQ4,
		   Q => NQ6
		   );
		 
U9 : registro  -- Registro de validaci�n
       port map (
		   ENTRADA => NQ6,
			SALIDA => NQ7,
			EN => NQ5,
			RCLK => CLK_OUT
			);
			
U10 : visualizacion   -- M�dulo de visualizaci�n
       port map (
		   E8 => NQ7(2 downto 0),
		   E7(0) => NQ7(28),
			E7(1) => NQ7(29),
			E7(2) => NQ7(30),
			E7(3) => '0',
			E6 => NQ7 (27 downto 24),       -- Desplazamos los datos con respecto a la                                            
			E5(0) => NQ7(21),               -- versi�n original
			E5(1) => NQ7(22),               -- de forma que los 14 primeros bits vayan
			E5(2) => NQ7(23),               -- al multiplexor 1
			E5(3) => '0',                   -- (correspondiente a la hora) y los 14 siguientes al 
			E4 => NQ7 (20 downto 17),       -- multiplexor 2 (correspondiente a la fecha)
		   E3(0) => NQ7(14),               -- los 3 �ltimos bits iran directamente al decodificador
			E3(1) => NQ7(15),               -- para ser decodificados y mandados a los LEDS de d�a de la semana
			E3(2) => NQ7(16),
			E3(3) => '0',
			E2 => NQ7 (13 downto 10),
			E1(0) => NQ7(7),
			E1(1) => NQ7(8),
			E1(2) => NQ7(9),
			E1(3) => '0',
			E0 => NQ7 (6 downto 3),
			PULSADOR => PULSADOR,
			CLK => CLK,
			LEDS => LEDS,
			SEG7 => SEG7,
			AN => AN
			);
			

end a_principal;